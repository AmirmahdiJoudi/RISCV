module controller ( 
    input [6:0] opcode, 
    input [2:0] func3,
    input [6:0] func7,

    input gt,
    input lt,
    input eq, 

    output PC_src,
    output jal_jalr,
    output alu_src1,
    output [1:0] alu_src2,
    output ensh2,
    output set0,
    output sgn_unsgn,
    output [2:0] imm_typ,
    output [3:0] alu_operation,
    output wb_src,
    output reg_write,
    output mem_read_i, 
    output mem_write_i,
    output b,
    output h,
    output w,
    output bhu,
    output IF_flush
);

    assign {IF_flush, PC_src, jal_jalr, alu_src1, alu_src2, ensh2, set0, sgn_unsgn, imm_typ, alu_operation, wb_src, reg_write, mem_read_i, mem_write_i, b, h, w, bhu} =
    // LUI
    (opcode==7'b0110111) ? 24'b0_0_0_0_01_0_0_0_100_0011_0_1_0_0_0_0_0_0 :
    // AUIPC
    (opcode==7'b0010111) ? 24'b0_0_0_1_01_0_0_0_100_0001_0_1_0_0_0_0_0_0 :
    // JAL
    (opcode==7'b1101111) ? 24'b1_1_0_1_10_0_0_0_101_0001_0_1_0_0_0_0_0_0 :
    // JALR
    (opcode==7'b1100111 && func3==3'b000) ? 24'b1_1_1_1_10_0_1_0_001_0001_0_1_0_0_0_0_0_0 :
    // BEQ
    (opcode==7'b1100011 && func3==3'b000) ? {eq, eq, 22'b0_0_00_0_0_0_011_0000_0_0_0_0_0_0_0_0} :
    // BNE
    (opcode==7'b1100011 && func3==3'b001) ? {~eq, ~eq, 22'b0_0_00_0_0_0_011_0000_0_0_0_0_0_0_0_0} :
    // BLT
    (opcode==7'b1100011 && func3==3'b100) ? {lt, lt, 22'b0_0_00_0_0_0_011_0000_0_0_0_0_0_0_0_0} :
    // BGE
    (opcode==7'b1100011 && func3==3'b101) ? {gt, gt, 22'b0_0_00_0_0_0_011_0000_0_0_0_0_0_0_0_0} :
    // BLTU
    (opcode==7'b1100011 && func3==3'b110) ? {lt, lt, 22'b0_0_00_0_0_1_011_0000_0_0_0_0_0_0_0_0} :
    // BGEU
    (opcode==7'b1100011 && func3==3'b111) ? {gt, gt, 22'b0_0_00_0_0_1_011_0000_0_0_0_0_0_0_0_0} :
    // LB
    (opcode==7'b0000011 && func3==3'b000) ? 24'b0_0_0_0_01_0_0_0_001_0001_1_1_1_0_1_0_0_0 :
    // LH
    (opcode==7'b0000011 && func3==3'b001) ? 24'b0_0_0_0_01_0_0_0_001_0001_1_1_1_0_0_1_0_0 :
    // LW
    (opcode==7'b0000011 && func3==3'b010) ? 24'b0_0_0_0_01_0_0_0_001_0001_1_1_1_0_0_0_1_0 :
    // LBU
    (opcode==7'b0000011 && func3==3'b100) ? 24'b0_0_0_0_01_0_0_0_001_0001_1_1_1_0_1_0_0_1 :
    // LHU
    (opcode==7'b0000011 && func3==3'b101) ? 24'b0_0_0_0_01_0_0_0_001_0001_1_1_1_0_0_1_0_1 :
    // SB
    (opcode==7'b0100011 && func3==3'b000) ? 24'b0_0_0_0_01_0_0_0_010_0001_0_0_0_1_1_0_0_0 :
    // SH
    (opcode==7'b0100011 && func3==3'b001) ? 24'b0_0_0_0_01_0_0_0_010_0001_0_0_0_1_0_1_0_0 :
    // SW
    (opcode==7'b0100011 && func3==3'b010) ? 24'b0_0_0_0_01_0_0_0_010_0001_0_0_0_1_0_0_1_0 :
    // ADDI
    (opcode==7'b0010011 && func3==3'b000) ? 24'b0_0_0_0_01_0_0_0_001_0001_0_1_0_0_0_0_0_0 :
    // SLTI
    (opcode==7'b0010011 && func3==3'b010) ? 24'b0_0_0_0_01_0_0_0_001_0100_0_1_0_0_0_0_0_0 :
    // SLTIU
    (opcode==7'b0010011 && func3==3'b011) ? 24'b0_0_0_0_01_0_0_0_001_0101_0_1_0_0_0_0_0_0 :
    // XORI
    (opcode==7'b0010011 && func3==3'b100) ? 24'b0_0_0_0_01_0_0_0_001_0110_0_1_0_0_0_0_0_0 :
    // ORI
    (opcode==7'b0010011 && func3==3'b110) ? 24'b0_0_0_0_01_0_0_0_001_0111_0_1_0_0_0_0_0_0 :
    // ANDI
    (opcode==7'b0010011 && func3==3'b111) ? 24'b0_0_0_0_01_0_0_0_001_1000_0_1_0_0_0_0_0_0 :
    // SLLI
    (opcode==7'b0010011 && func3==3'b001 && func7==7'b0000000) ? 24'b0_0_0_0_01_0_0_0_110_1001_0_1_0_0_0_0_0_0 :
    // SRLI
    (opcode==7'b0010011 && func3==3'b101 && func7==7'b0000000) ? 24'b0_0_0_0_01_0_0_0_110_1010_0_1_0_0_0_0_0_0 :
    // SRAI
    (opcode==7'b0010011 && func3==3'b101 && func7==7'b0100000) ? 24'b0_0_0_0_01_0_0_0_110_1011_0_1_0_0_0_0_0_0 :
    // ADD
    (opcode==7'b0110011 && func3==3'b000 && func7==7'b0000000) ? 24'b0_0_0_0_00_0_0_0_000_0001_0_1_0_0_0_0_0_0 :
    // SUB
    (opcode==7'b0110011 && func3==3'b000 && func7==7'b0100000) ? 24'b0_0_0_0_00_0_0_0_000_0010_0_1_0_0_0_0_0_0 :
    // SLL
    (opcode==7'b0110011 && func3==3'b001 && func7==7'b0000000) ? 24'b0_0_0_0_00_0_0_0_000_1001_0_1_0_0_0_0_0_0 :
    // SLT
    (opcode==7'b0110011 && func3==3'b010 && func7==7'b0000000) ? 24'b0_0_0_0_00_0_0_0_000_0100_0_1_0_0_0_0_0_0 :
    // SLTU
    (opcode==7'b0110011 && func3==3'b011 && func7==7'b0000000) ? 24'b0_0_0_0_00_0_0_0_000_0101_0_1_0_0_0_0_0_0 :
    // XOR
    (opcode==7'b0110011 && func3==3'b100 && func7==7'b0000000) ? 24'b0_0_0_0_00_0_0_0_000_0110_0_1_0_0_0_0_0_0 :
    // SRL
    (opcode==7'b0110011 && func3==3'b101 && func7==7'b0000000) ? 24'b0_0_0_0_00_0_0_0_000_1010_0_1_0_0_0_0_0_0 :
    // SRA
    (opcode==7'b0110011 && func3==3'b101 && func7==7'b0100000) ? 24'b0_0_0_0_00_0_0_0_000_1011_0_1_0_0_0_0_0_0 :
    // OR
    (opcode==7'b0110011 && func3==3'b110 && func7==7'b0000000) ? 24'b0_0_0_0_00_0_0_0_000_0111_0_1_0_0_0_0_0_0 :
    // AND
    (opcode==7'b0110011 && func3==3'b111 && func7==7'b0000000) ? 24'b0_0_0_0_00_0_0_0_000_1000_0_1_0_0_0_0_0_0 :
    
    24'b0_0_0_0_00_0_0_0_000_0000_0_0_0_0_0_0_0_0;

endmodule
